module bcd_conv(c0,s3,s2,s1,s0,z2,y2,x2,w2,z1,y1,x1,w1);
input c0,s3,s2,s1,s0;
output z2,x2,y2,w2,z1,x1,y1,w1;
reg z2,x2,y2,w2,z1,x1,y1,w1;

always@(z2 or y2 or w2 or z1 or y1 or x1 or w1)
 case ({c0,s3,s2,s1,s0})
  5'b00000:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00000000;
  5'b00001:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00000001;
  5'b00010:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00000010;
  5'b00011:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00000011;
  5'b00100:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00000100;
  5'b00101:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00000101;
  5'b00110:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00000110;
  5'b00111:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00000111;
  5'b01000:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00001000;
  5'b01001:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00001001;
  5'b01010:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00010000;
  5'b01011:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00010001;
  5'b01100:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00010010;
  5'b01101:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00010011;
  5'b01110:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00010100;
  5'b01111:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00010101;
  5'b10000:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00010110;
  5'b10001:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00010111;
  5'b10010:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00011000;
  5'b10011:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00011001;
  5'b10100:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00100000;
  5'b10101:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00100001;
  5'b10110:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00100010;
  5'b10111:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00100011;
  5'b11000:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00100100;
  5'b11001:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00100101;
  5'b11010:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00100110;
  5'b11011:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00100111;
  5'b11100:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00101000;
  5'b11101:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00101001;
  5'b11110:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00110000;
  5'b11111:{z2,y2,x2,w2,z1,y1,x1,w1} = 8'b00110001;
  endcase
  
  endmodule