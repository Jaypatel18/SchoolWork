module Decoder16bit (WA, WR, R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15);
	input [3:0] WA; 
	input WR;
	output R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15;
	reg R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15;
	
	always@(WA[3] or WA[2] or WA[1] or WA[0] or WR)
	begin
		case({WR, WA[3], WA[2], WA[1], WA[0]})
			5'b00000:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000000000;
			5'b00001:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000000000;
			5'b00010:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000000000;
			5'b00011:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000000000;
			5'b00100:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000000000;
			5'b00101:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000000000;
			5'b00110:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000000000;
			5'b00111:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000000000;
			5'b01000:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000000000;
			5'b01001:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000000000;
			5'b01010:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000000000;
			5'b01011:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000000000;
			5'b01100:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000000000;
			5'b01101:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000000000;
			5'b01110:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000000000;
			5'b01111:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000000000;
			5'b10000:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b1000000000000000;
			5'b10001:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0100000000000000;
			5'b10010:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0010000000000000;
			5'b10011:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0001000000000000;
			5'b10100:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000100000000000;
			5'b10101:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000010000000000;
			5'b10110:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000001000000000;
			5'b10111:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000100000000;
			5'b11000:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000010000000;
			5'b11001:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000001000000;
			5'b11010:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000100000;
			5'b11011:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000010000;
			5'b11100:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000001000;
			5'b11101:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000000100;
			5'b11110:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000000010;
			5'b11111:{R00, R01, R02, R03, R04, R05, R06, R07, R08, R09, R10, R11, R12, R13, R14, R15}=16'b0000000000000001;
		endcase
	end
	
endmodule